`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Design Name: 
// Module Name: fbe_pkg
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////
//package fbe_pkg;

    parameter ECHO_AND_INIT_COEFF = 9;
    parameter ECHO_IN_GAIN_FDB_GAIN = 13;
    parameter FDB_DELAY_FB_GAIN = 17;
    parameter LP_ORDER_GAIN = 21;
    parameter BP_ORDER_GAIN = 25;
    parameter HP_ORDER_GAIN = 29;
    
//endpackage
